//UNSIGNED MULTIPLIER
module multiplier (multiplier, multiplicand, product);
  parameter parallelism=8;
  parameter ARCH_TYPE=0;
  /*SELECT ARCH_TYPE IN MOSULE INSTANCE AS:
      0 : synthesizer choose
      1 : complete csa implmentation
      2 : row cutted implmentation*/

  input signed [parallelism-1:0] multiplier;
  input signed [parallelism-1:0] multiplicand;
  output signed [2*parallelism-1:0] product;
  
  //needed for Sign&Magnitude multiplier
  logic sign;
  logic unsigned [parallelism-2:0] SM_multiplier;
  logic unsigned [parallelism-2:0] SM_multiplicand;
  logic unsigned [2*(parallelism-1)-1:0] SM_product;
  logic unsigned [2*(parallelism-1)-1:0] r_prod; //last parallelism-2 lenght of product
  
  //needed for csaTree
  logic signed [parallelism-1:0] pps    [parallelism-1:0];
  logic signed [parallelism*2-1:0] sums   [parallelism-2:0];
  logic signed [parallelism*2-1:0] carrys [parallelism-2:0];

  genvar i;
  generate
    if (ARCH_TYPE==0) begin: beha //synthesizer choose
      assign product = multiplier*multiplicand;
    end
    else if (ARCH_TYPE==1) begin: csaHandWritten //complete csa tree
      //generate partial products
      for (i=0;i<parallelism;i++) begin
        assign pps[i] = (multiplier[i]) ? multiplicand : 8'b0;
      end
      //building the tree
      assign product[0] = pps[0][0];
      csaRow #(parallelism-1) row1 (  .a(pps[0][parallelism-1:1]),
                                      .b(pps[1][parallelism-2:0]),
                                      .ci(7'b0),
                                      .s({sums[0],product[1]}),
                                      .co(carrys[0]));
      //make all the following lines exept for last carry adder!
      for (i=1;i<parallelism-1;i++) begin
        csaRow #(parallelism-1) row1 (  .a(pps[i+1][parallelism-2:0]),
                                        .b({pps[i][parallelism-1],sums[i-1][parallelism-3:0]}),
                                        .ci(carrys[i-1][parallelism-2:0]),
                                        .s({sums[i],product[i+1]}),
                                        .co(carrys[i]));
      end
      //adder for last row
      adder #(.parallelism(parallelism),
              .ARCH_TYPE(1)) rcaFinale (.add1({1'b0,pps[parallelism-1][parallelism-1],sums[parallelism-2]}),
                                        .add0({1'b0,carrys[parallelism-2]}),
                                        .carry_in(1'b0),
                                        .sum(product[2*parallelism-1:parallelism]));
    end
    else if (ARCH_TYPE==2) begin: csaAuto //autogenerated arhitecture
      //generate partial products
      for (i=0;i<parallelism;i++) begin
        assign pps[i] = (multiplier[i]) ? multiplicand : 8'b0;
      end
      //AUTO_PRINT
    end
    else if (ARCH_TYPE==3) begin: behaSM //behavioural Sing and magnitude
      // NOTE that in such implementation multiplier and multiplicand are already given in S&M format
      assign SM_multiplicand = multiplicand[parallelism-2:0];
      assign SM_multiplier = multiplier[parallelism-2:0];
      assign SM_product = SM_multiplier*SM_multiplicand;
      assign sign = multiplicand[parallelism-1] ^ multiplier[parallelism-1];
      assign product [2*parallelism -1:2*parallelism -2] = {2{sign}}; //sign for the first two bit of product
      assign r_prod = SM_product^{ $size(SM_product){sign}};
      assign product [2*parallelism - 3:0] = r_prod;
    end
  endgenerate
endmodule //multiplier
