//UNSIGNED MULTIPLIER
module multiplier (multiplier, multiplicand, product);
  parameter parallelism=8;
  parameter ARCH_TYPE=0;
  /*SELECT ARCH_TYPE IN MOSULE INSTANCE AS:
      0 : synthesizer choose
      1 : complete csa implmentation
      2 : row cutted implmentation*/

  input unsigned [parallelism-1:0] multiplier;
  input unsigned [parallelism-1:0] multiplicand;
  output unsigned [2*parallelism-1:0] product;

  logic unsigned [parallelism-1:0] pps    [parallelism-1:0];
  logic unsigned [parallelism*2-1:0] sums   [parallelism-2:0];
  logic unsigned [parallelism*2-1:0] carrys [parallelism-2:0];

  genvar i;
  generate
    if (ARCH_TYPE==0) begin: beha //synthesizer choose
      assign product = multiplier*multiplicand;
    end
    else if (ARCH_TYPE==1) begin: csaHandWritten //complete csa tree
      //generate partial products
      for (i=0;i<parallelism;i++) begin
        assign pps[i] = (multiplier[i]) ? multiplicand : 8'b0;
      end
      //building the tree
      assign product[0] = pps[0][0];
      csaRow #(parallelism-1) row1 (  .a(pps[0][parallelism-1:1]),
                                      .b(pps[1][parallelism-2:0]),
                                      .ci(7'b0),
                                      .s({sums[0],product[1]}),
                                      .co(carrys[0]));
      //make all the following lines exept for last carry adder!
      for (i=1;i<parallelism-1;i++) begin
        csaRow #(parallelism-1) row1 (  .a(pps[i+1][parallelism-2:0]),
                                        .b({pps[i][parallelism-1],sums[i-1][parallelism-3:0]}),
                                        .ci(carrys[i-1][parallelism-2:0]),
                                        .s({sums[i],product[i+1]}),
                                        .co(carrys[i]));
      end
      //adder for last row
      adder #(.parallelism(parallelism),
              .ARCH_TYPE(1)) rcaFinale (.add1({1'b0,pps[parallelism-1][parallelism-1],sums[parallelism-2]}),
                                        .add0({1'b0,carrys[parallelism-2]}),
                                        .carry_in(1'b0),
                                        .sum(product[2*parallelism-1:parallelism]));
    end
    else if (ARCH_TYPE==2) begin: csaAuto //autogenerated arhitecture
      //generate partial products
      for (i=0;i<parallelism;i++) begin
        assign pps[i] = (multiplier[i]) ? multiplicand : 8'b0;
      end
assign product[0] = 1'b0;
assign product[1] = pps[1][0];
fullAdder fh0 (.a(pps[1][1]),.b(pps[2][0]),.ci(1'b0),.s(sums[0][0]),.co(carrys[0][0]));
fullAdder fh1 (.a(pps[1][2]),.b(pps[2][1]),.ci(1'b0),.s(sums[0][1]),.co(carrys[0][1]));
fullAdder fh2 (.a(pps[1][3]),.b(pps[2][2]),.ci(pps[4][0]),.s(sums[0][2]),.co(carrys[0][2]));
fullAdder fh3 (.a(pps[1][4]),.b(pps[2][3]),.ci(pps[4][1]),.s(sums[0][3]),.co(carrys[0][3]));
fullAdder fh4 (.a(pps[1][5]),.b(pps[2][4]),.ci(pps[4][2]),.s(sums[0][4]),.co(carrys[0][4]));
fullAdder fh5 (.a(pps[1][6]),.b(pps[2][5]),.ci(pps[4][3]),.s(sums[0][5]),.co(carrys[0][5]));
fullAdder fh6 (.a(pps[1][7]),.b(pps[2][6]),.ci(pps[4][4]),.s(sums[0][6]),.co(carrys[0][6]));
fullAdder fh7 (.a(1'b0),.b(pps[2][7]),.ci(pps[4][5]),.s(sums[0][7]),.co(carrys[0][7]));
fullAdder fh8 (.a(1'b0),.b(1'b0),.ci(pps[4][6]),.s(sums[0][8]),.co(carrys[0][8]));
fullAdder fh9 (.a(1'b0),.b(1'b0),.ci(pps[4][7]),.s(sums[0][9]),.co(carrys[0][9]));
assign product[2] = sums[0][0];
fullAdder fh10 (.a(sums[0][1]),.b(carrys[0][0]),.ci(1'b0),.s(sums[1][0]),.co(carrys[1][0]));
fullAdder fh11 (.a(sums[0][2]),.b(carrys[0][1]),.ci(1'b0),.s(sums[1][1]),.co(carrys[1][1]));
fullAdder fh12 (.a(sums[0][3]),.b(carrys[0][2]),.ci(pps[5][0]),.s(sums[1][2]),.co(carrys[1][2]));
fullAdder fh13 (.a(sums[0][4]),.b(carrys[0][3]),.ci(pps[5][1]),.s(sums[1][3]),.co(carrys[1][3]));
fullAdder fh14 (.a(sums[0][5]),.b(carrys[0][4]),.ci(pps[5][2]),.s(sums[1][4]),.co(carrys[1][4]));
fullAdder fh15 (.a(sums[0][6]),.b(carrys[0][5]),.ci(pps[5][3]),.s(sums[1][5]),.co(carrys[1][5]));
fullAdder fh16 (.a(sums[0][7]),.b(carrys[0][6]),.ci(pps[5][4]),.s(sums[1][6]),.co(carrys[1][6]));
fullAdder fh17 (.a(sums[0][8]),.b(carrys[0][7]),.ci(pps[5][5]),.s(sums[1][7]),.co(carrys[1][7]));
fullAdder fh18 (.a(sums[0][9]),.b(carrys[0][8]),.ci(pps[5][6]),.s(sums[1][8]),.co(carrys[1][8]));
fullAdder fh19 (.a(1'b0),.b(carrys[0][9]),.ci(pps[5][7]),.s(sums[1][9]),.co(carrys[1][9]));
assign product[3] = sums[1][0];
fullAdder fh20 (.a(sums[1][1]),.b(carrys[1][0]),.ci(1'b0),.s(sums[2][0]),.co(carrys[2][0]));
fullAdder fh21 (.a(sums[1][2]),.b(carrys[1][1]),.ci(1'b0),.s(sums[2][1]),.co(carrys[2][1]));
fullAdder fh22 (.a(sums[1][3]),.b(carrys[1][2]),.ci(pps[6][0]),.s(sums[2][2]),.co(carrys[2][2]));
fullAdder fh23 (.a(sums[1][4]),.b(carrys[1][3]),.ci(pps[6][1]),.s(sums[2][3]),.co(carrys[2][3]));
fullAdder fh24 (.a(sums[1][5]),.b(carrys[1][4]),.ci(pps[6][2]),.s(sums[2][4]),.co(carrys[2][4]));
fullAdder fh25 (.a(sums[1][6]),.b(carrys[1][5]),.ci(pps[6][3]),.s(sums[2][5]),.co(carrys[2][5]));
fullAdder fh26 (.a(sums[1][7]),.b(carrys[1][6]),.ci(pps[6][4]),.s(sums[2][6]),.co(carrys[2][6]));
fullAdder fh27 (.a(sums[1][8]),.b(carrys[1][7]),.ci(pps[6][5]),.s(sums[2][7]),.co(carrys[2][7]));
fullAdder fh28 (.a(sums[1][9]),.b(carrys[1][8]),.ci(pps[6][6]),.s(sums[2][8]),.co(carrys[2][8]));
fullAdder fh29 (.a(1'b0),.b(carrys[1][9]),.ci(pps[6][7]),.s(sums[2][9]),.co(carrys[2][9]));
assign product[4] = sums[2][0];
fullAdder fh30 (.a(sums[2][1]),.b(carrys[2][0]),.ci(1'b0),.s(sums[3][0]),.co(carrys[3][0]));
fullAdder fh31 (.a(sums[2][2]),.b(carrys[2][1]),.ci(1'b0),.s(sums[3][1]),.co(carrys[3][1]));
fullAdder fh32 (.a(sums[2][3]),.b(carrys[2][2]),.ci(pps[7][0]),.s(sums[3][2]),.co(carrys[3][2]));
fullAdder fh33 (.a(sums[2][4]),.b(carrys[2][3]),.ci(pps[7][1]),.s(sums[3][3]),.co(carrys[3][3]));
fullAdder fh34 (.a(sums[2][5]),.b(carrys[2][4]),.ci(pps[7][2]),.s(sums[3][4]),.co(carrys[3][4]));
fullAdder fh35 (.a(sums[2][6]),.b(carrys[2][5]),.ci(pps[7][3]),.s(sums[3][5]),.co(carrys[3][5]));
fullAdder fh36 (.a(sums[2][7]),.b(carrys[2][6]),.ci(pps[7][4]),.s(sums[3][6]),.co(carrys[3][6]));
fullAdder fh37 (.a(sums[2][8]),.b(carrys[2][7]),.ci(pps[7][5]),.s(sums[3][7]),.co(carrys[3][7]));
fullAdder fh38 (.a(sums[2][9]),.b(carrys[2][8]),.ci(pps[7][6]),.s(sums[3][8]),.co(carrys[3][8]));
fullAdder fh39 (.a(1'b0),.b(carrys[2][9]),.ci(pps[7][7]),.s(sums[3][9]),.co(carrys[3][9]));
assign product[5] = sums[3][0];
adder #(.parallelism(10),.ARCH_TYPE(1)) adder (.add1({1'b0,sums[3][9:1]}),.add0(carrys[3][9:0]),.carry_in(1'b0),.sum(product[15:6]));
    end
  endgenerate
endmodule //multiplier
